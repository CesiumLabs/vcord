module valkyria

pub struct Ready {
pub mut:
        v          int
        session_id string
        shard      []int
}